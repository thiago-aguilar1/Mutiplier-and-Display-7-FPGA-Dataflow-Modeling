module multiplicador (
						input [4:0] A,   // tem 5 bits
						output a1, b1, c1, d1, e1, f1, g1, a2, b2, c2, d2, e2, f2, g2, 
							   a3, b3, c3, d3, e3, f3, g3, a4, b4, c4, d4, e4, f4, g4 
						);
						   //o valor m�ximo de A � 31, e 31*3=93 , logo,
						   //o produto m�ximo tamb�m poder� ser mostrado nos displays.
wire [6:0]  seteSegmentos1,		
			seteSegmentos2,
			seteSegmentos3,
			seteSegmentos4;				


assign {seteSegmentos2, seteSegmentos1} = (A == 5'b00_000) ? {7'b1111_110, 7'b1111_110} :  //0
										  (A == 5'b00_001) ? {7'b1111_110, 7'b0110_000} :  //1
										  (A == 5'b00_010) ? {7'b1111_110, 7'b1101_101} :  //2
										  (A == 5'b00_011) ? {7'b1111_110, 7'b1111_001} :  //3
										  (A == 5'b00_100) ? {7'b1111_110, 7'b0110_011} :  //4
										  (A == 5'b00_101) ? {7'b1111_110, 7'b1011_011} :  //5
										  (A == 5'b00_110) ? {7'b1111_110, 7'b1011_111} :  //6
										  (A == 5'b00_111) ? {7'b1111_110, 7'b1110_000} :  //7
										  (A == 5'b01_000) ? {7'b1111_110, 7'b1111_111} :  //8
										  (A == 5'b01_001) ? {7'b1111_110, 7'b1111_011} :  //9
										  (A == 5'b01_010) ? {7'b0110_000, 7'b1111_110} :  //10
										  (A == 5'b01_011) ? {7'b0110_000, 7'b0110_000} :  //11
										  (A == 5'b01_100) ? {7'b0110_000, 7'b1101_101} :  //12
										  (A == 5'b01_101) ? {7'b0110_000, 7'b1111_001} :  //13
										  (A == 5'b01_110) ? {7'b0110_000, 7'b0110_011} :  //14
										  (A == 5'b01_111) ? {7'b0110_000, 7'b1011_011} :  //15
										  (A == 5'b10_000) ? {7'b0110_000, 7'b1011_111} :  //16
										  (A == 5'b10_001) ? {7'b0110_000, 7'b1110_000} :  //17
										  (A == 5'b10_010) ? {7'b0110_000, 7'b1111_111} :  //18
										  (A == 5'b10_011) ? {7'b0110_000, 7'b1111_011} :  //19
										  (A == 5'b10_100) ? {7'b1101_101, 7'b1111_110} :  //20
										  (A == 5'b10_101) ? {7'b1101_101, 7'b0110_000} :  //21
										  (A == 5'b10_110) ? {7'b1101_101, 7'b1101_101} :  //22
										  (A == 5'b10_111) ? {7'b1101_101, 7'b1111_001} :  //23
										  (A == 5'b11_000) ? {7'b1101_101, 7'b0110_011} :  //24
										  (A == 5'b11_001) ? {7'b1101_101, 7'b1011_011} :  //25
										  (A == 5'b11_010) ? {7'b1101_101, 7'b1011_111} :  //26
										  (A == 5'b11_011) ? {7'b1101_101, 7'b1110_000} :  //27
										  (A == 5'b11_100) ? {7'b1101_101, 7'b1111_111} :  //28
										  (A == 5'b11_101) ? {7'b1101_101, 7'b1111_011} :  //29
										  (A == 5'b11_110) ? {7'b1111_001, 7'b1111_110} :  //30
										  (A == 5'b11_111) ? {7'b1111_001, 7'b0110_000} :  //31
										  {7'b0000_000, 7'b0000_000};  
										  
										  

assign {a2, b2, c2, d2, e2, f2, g2, a1, b1, c1, d1, e1, f1, g1} = {seteSegmentos2, seteSegmentos1};



assign {seteSegmentos4, seteSegmentos3} = (A == 5'b00_000) ? {7'b1111_110, 7'b1111_110} :  //0
										  (A == 5'b00_001) ? {7'b1111_110, 7'b1111_001} :  //3
										  (A == 5'b00_010) ? {7'b1111_110, 7'b1011_111} :  //6
										  (A == 5'b00_011) ? {7'b1111_110, 7'b1111_011} :  //9
										  (A == 5'b00_100) ? {7'b0110_000, 7'b1101_101} :  //12
										  (A == 5'b00_101) ? {7'b0110_000, 7'b1011_011} :  //15
										  (A == 5'b00_110) ? {7'b0110_000, 7'b1111_111} :  //18
										  (A == 5'b00_111) ? {7'b1101_101, 7'b0110_000} :  //21
										  (A == 5'b01_000) ? {7'b1101_101, 7'b0110_011} :  //24
										  (A == 5'b01_001) ? {7'b1101_101, 7'b1110_000} :  //27
										  (A == 5'b01_010) ? {7'b1111_001, 7'b1111_110} :  //30
										  (A == 5'b01_011) ? {7'b1111_001, 7'b1111_001} :  //33
										  (A == 5'b01_100) ? {7'b1111_001, 7'b1011_111} :  //36
										  (A == 5'b01_101) ? {7'b1111_001, 7'b1111_011} :  //39
										  (A == 5'b01_110) ? {7'b0110_011, 7'b1101_101} :  //42
										  (A == 5'b01_111) ? {7'b0110_011, 7'b1011_011} :  //45
										  (A == 5'b10_000) ? {7'b0110_011, 7'b1111_111} :  //48
										  (A == 5'b10_001) ? {7'b1011_011, 7'b0110_000} :  //51
										  (A == 5'b10_010) ? {7'b1011_011, 7'b0110_011} :  //54
										  (A == 5'b10_011) ? {7'b1011_011, 7'b1110_000} :  //57
										  (A == 5'b10_100) ? {7'b1011_111, 7'b1111_110} :  //60
										  (A == 5'b10_101) ? {7'b1011_111, 7'b1111_001} :  //63
										  (A == 5'b10_110) ? {7'b1011_111, 7'b1011_111} :  //66
										  (A == 5'b10_111) ? {7'b1011_111, 7'b1111_011} :  //69
										  (A == 5'b11_000) ? {7'b1110_000, 7'b1101_101} :  //72
										  (A == 5'b11_001) ? {7'b1110_000, 7'b1011_011} :  //75
										  (A == 5'b11_010) ? {7'b1110_000, 7'b1111_111} :  //78
										  (A == 5'b11_011) ? {7'b1111_111, 7'b0110_000} :  //81
										  (A == 5'b11_100) ? {7'b1111_111, 7'b0110_011} :  //84
										  (A == 5'b11_101) ? {7'b1111_111, 7'b1110_000} :  //87
										  (A == 5'b11_110) ? {7'b1111_011, 7'b1111_110} :  //90
										  (A == 5'b11_111) ? {7'b1111_011, 7'b1111_001} :  //93
										  {7'b0000_000, 7'b0000_000};  
										  
										  

assign {a4, b4, c4, d4, e4, f4, g4, a3, b3, c3, d3, e3, f3, g3} = {seteSegmentos4, seteSegmentos3};

endmodule   

